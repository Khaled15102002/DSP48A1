module DSP(A, B, C, D, CARRYIN, M, P, CARRYOUT, CARRYOUTF, CLK, OPMODE, BCIN, 
CEA, CEB, CEC, CECARRYIN, CED, CEM, CEOPMODE, CEP, RSTA, RSTB, RSTC, RSTCARRYIN, RSTD, RSTM, RSTOPMODE, RSTP, BCOUT, PCIN, PCOUT); 
localparam SYNC = 0, ASYNC = 1, OPMODE5 = 0, CARRYIn = 1, CASCODE = 1, DIRECT = 0;
parameter A0REG = 0, A1REG = 1, B0REG = 0, B1REG = 1;
parameter CREG = 1, DREG = 1, MREG = 1, PREG = 1, CARRYINREG = 1, CARRYOUTREG = 1, OPMODEREG = 1;
parameter CARRYINSEL = OPMODE5;
parameter B_INPUT = DIRECT;
parameter RSTTYPE = SYNC;
parameter A_WIDTH = 18, B_WIDTH = 18, C_WIDTH = 48, D_WIDTH = 18, M_WIDTH = 36, P_WIDTH = 48, OPMODE_WIDTH = 8;
input [17:0] A, B, BCIN;
input [17:0] D;
input [47:0] C, PCIN;
input CARRYIN, CLK, CEA, CEB, CEC, CECARRYIN, CED, CEM, CEOPMODE, CEP;
input RSTA, RSTB, RSTC, RSTCARRYIN, RSTD, RSTM, RSTOPMODE, RSTP;
input [7:0] OPMODE;
output [35:0] M;
output [47:0] P, PCOUT;
output CARRYOUT, CARRYOUTF;
output [17:0] BCOUT;
wire [7:0] OPMODE_out;
wire [17:0] A_mux_out, B_mux_out, MUX0B_out;
wire [17:0] D_mux_out;
wire [47:0] C_mux_out, X_mux_out, Z_mux_out, PRE_ADDER_SUB_2;
wire [17:0] PRE_ADDER_SUB_1, MUX_OP4, MULTI_1, MULTI_2;
wire [35:0] MULTI;
wire [47:0] M_ex;
wire Carry_Cascode_in, CIN, Carry_Cascode_out;
REG_MUX #(OPMODE_WIDTH,RSTTYPE,OPMODEREG) x0 (OPMODE, CLK, RSTOPMODE, CEOPMODE, OPMODE_out);
REG_MUX #(D_WIDTH,RSTTYPE,DREG) x1 (D, CLK, RSTD, CED, D_mux_out);
REG_MUX #(A_WIDTH,RSTTYPE,A0REG) x2 (A, CLK, RSTA, CEA, A_mux_out);
REG_MUX #(C_WIDTH,RSTTYPE,CREG) x3 (C, CLK, RSTC, CEC, C_mux_out);
assign MUX0B_out = (B_INPUT == DIRECT)? B : (B_INPUT == CASCODE)? BCIN : 0;
REG_MUX #(B_WIDTH,RSTTYPE,B0REG) x5 (MUX0B_out, CLK, RSTB, CEB, B_mux_out);
assign PRE_ADDER_SUB_1 = (OPMODE_out[6])? D_mux_out-B_mux_out : D_mux_out+B_mux_out;
assign MUX_OP4 = (OPMODE_out[4])? PRE_ADDER_SUB_1 : B_mux_out;
REG_MUX #(B_WIDTH,RSTTYPE,B1REG) x6 (MUX_OP4, CLK, RSTB, CEB, MULTI_1);
REG_MUX #(A_WIDTH,RSTTYPE,A1REG) x7 (A_mux_out, CLK, RSTA, CEA, MULTI_2);
assign BCOUT = MULTI_1;
assign MULTI = MULTI_1 * MULTI_2;
REG_MUX #(M_WIDTH,RSTTYPE,MREG) x8 (MULTI, CLK, RSTM, CEM, M);
assign Carry_Cascode_in = (CARRYINSEL==OPMODE5)? OPMODE_out[5] : (CARRYINSEL==CARRYIn)? CARRYIN : 0;
REG_MUX #(1,RSTTYPE,CARRYINREG) x9 (Carry_Cascode_in, CLK, RSTCARRYIN, CECARRYIN, CIN);
assign M_ex = {{12{1'b0}},M};
assign X_mux_out = (OPMODE_out[1:0]==3)? {D[11:0],A,B} : (OPMODE_out[1:0]==2)? P : (OPMODE_out[1:0]==1)? M_ex : 0;
assign Z_mux_out = (OPMODE_out[3:2]==3)? C_mux_out : (OPMODE_out[3:2]==2)? P : (OPMODE_out[3:2]==1)? PCIN : 0;
assign {Carry_Cascode_out,PRE_ADDER_SUB_2} = (OPMODE_out[7]==0)? (X_mux_out + Z_mux_out + CIN) : (Z_mux_out-(X_mux_out+CIN));
REG_MUX #(1,RSTTYPE,CARRYOUTREG) x10 (Carry_Cascode_out, CLK, RSTCARRYIN, CECARRYIN, CARRYOUT);
REG_MUX #(P_WIDTH,RSTTYPE,PREG) x11 (PRE_ADDER_SUB_2, CLK, RSTP, CEP, P);
assign CARRYOUTF = CARRYOUT;
assign PCOUT = P;
endmodule

